library verilog;
use verilog.vl_types.all;
entity menorq_vlg_vec_tst is
end menorq_vlg_vec_tst;

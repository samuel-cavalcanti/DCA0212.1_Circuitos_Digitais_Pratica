library verilog;
use verilog.vl_types.all;
entity memoria_de_instrucoes_vlg_vec_tst is
end memoria_de_instrucoes_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity unidade_de_controle_vlg_vec_tst is
end unidade_de_controle_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity mux_3x1_vlg_vec_tst is
end mux_3x1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ffd_vlg_vec_tst is
end ffd_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity inverter_vlg_vec_tst is
end inverter_vlg_vec_tst;

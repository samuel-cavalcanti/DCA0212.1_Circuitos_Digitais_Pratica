library verilog;
use verilog.vl_types.all;
entity somador_complemento_de_2_vlg_vec_tst is
end somador_complemento_de_2_vlg_vec_tst;

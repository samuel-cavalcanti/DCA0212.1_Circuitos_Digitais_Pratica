library verilog;
use verilog.vl_types.all;
entity decision_controller_vlg_vec_tst is
end decision_controller_vlg_vec_tst;

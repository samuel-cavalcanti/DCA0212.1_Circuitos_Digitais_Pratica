library verilog;
use verilog.vl_types.all;
entity contraction_vlg_vec_tst is
end contraction_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity bloco_operacional_vlg_vec_tst is
end bloco_operacional_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity decodificador_vlg_vec_tst is
end decodificador_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity banco_de_registradores_vlg_vec_tst is
end banco_de_registradores_vlg_vec_tst;

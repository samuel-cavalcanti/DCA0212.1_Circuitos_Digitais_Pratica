library verilog;
use verilog.vl_types.all;
entity pacemaker_vlg_vec_tst is
end pacemaker_vlg_vec_tst;

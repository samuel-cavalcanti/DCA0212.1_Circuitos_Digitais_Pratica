library ieee;
use ieee.std_logic_1164.all; 


entity display is 
port ( distance : in std_logic_vector (8 downto 0);
		 thousands_display: out std_logic_vector(6 downto 0 ); -- hex3
		 hundreds_display : out std_logic_vector(6 downto 0 ); -- hex2
		 tens_display : out std_logic_vector(6 downto 0 ); -- hex1
		 units_display : out std_logic_vector(6 downto 0 )); -- hex0
		  
end entity;


architecture behavior of display is 

type decimal_places_type is array(0 to 3) of std_logic_vector(3 downto 0);
type display_places_type is array(0 to 3) of std_logic_vector(6 downto 0 );

signal decimal_places : decimal_places_type;
signal display_places : display_places_type;



begin

 binary_to_decimal : entity work.binary_to_decimal(behavior)
								port map ( distance=>distance,
											  units_mm => decimal_places(0),
											  tens_mm => decimal_places(1),
											  hundreds_mm => decimal_places(2),
											  thousands_mm => decimal_places(3));

 seven_segments_generate: for i in 0 to 3 generate
					seven_segments: entity work.decodificador(table)
							port map(s => decimal_places(i),
										h => display_places(i));
					end generate seven_segments_generate;
										
units_display<= display_places(0);
tens_display <= display_places(1);
hundreds_display <= display_places(2);
thousands_display <= display_places(3);




end architecture;
library verilog;
use verilog.vl_types.all;
entity utrassonic_sensor_vlg_vec_tst is
end utrassonic_sensor_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity bloco_de_controle_vlg_vec_tst is
end bloco_de_controle_vlg_vec_tst;

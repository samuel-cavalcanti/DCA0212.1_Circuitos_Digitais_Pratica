library verilog;
use verilog.vl_types.all;
entity contador_de_programa_vlg_vec_tst is
end contador_de_programa_vlg_vec_tst;

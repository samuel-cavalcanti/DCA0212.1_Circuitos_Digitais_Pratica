library verilog;
use verilog.vl_types.all;
entity button_vlg_sample_tst is
    port(
        key_0           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end button_vlg_sample_tst;

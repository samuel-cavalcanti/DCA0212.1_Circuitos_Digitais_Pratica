library verilog;
use verilog.vl_types.all;
entity registrador_de_instrucao_vlg_vec_tst is
end registrador_de_instrucao_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity button_vlg_vec_tst is
end button_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity memoriaD_vlg_vec_tst is
end memoriaD_vlg_vec_tst;

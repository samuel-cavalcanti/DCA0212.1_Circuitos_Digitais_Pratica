library verilog;
use verilog.vl_types.all;
entity maiorq_vlg_check_tst is
    port(
        resultmaq       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end maiorq_vlg_check_tst;

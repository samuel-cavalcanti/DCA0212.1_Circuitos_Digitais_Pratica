library verilog;
use verilog.vl_types.all;
entity contraction_vlg_check_tst is
    port(
        p               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end contraction_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity processador_programavel_vlg_vec_tst is
end processador_programavel_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity processador_programavel_vlg_sample_tst is
    port(
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end processador_programavel_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity menorq_vlg_check_tst is
    port(
        resultmeq       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end menorq_vlg_check_tst;

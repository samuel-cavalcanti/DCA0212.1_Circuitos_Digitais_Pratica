library verilog;
use verilog.vl_types.all;
entity maiorq_vlg_vec_tst is
end maiorq_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity set_clock_vlg_vec_tst is
end set_clock_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity trigger_control_vlg_vec_tst is
end trigger_control_vlg_vec_tst;

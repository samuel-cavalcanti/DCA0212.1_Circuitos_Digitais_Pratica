library verilog;
use verilog.vl_types.all;
entity comparador_vlg_vec_tst is
end comparador_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity button_vlg_check_tst is
    port(
        keyonoff        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end button_vlg_check_tst;
